module(input bit[31:0] inp_reg1,
	input bit[31:0] inp_reg2,
	output logic bit[31:0] out_reg);
	
endmodule
